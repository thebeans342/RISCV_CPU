module PC_reg (
    input logic 
)