module ALU (
    input logic op1,
    input logic op2,
    input logic ALUctrl,
    output logic ALUout,
    output logic EQ
)
